
`include "../env/svbt_interface.sv"
`include "../env/svbt_base_unit.sv"
`include "../env/svbt_packet.sv"
`include "../env/svbt_reset_bfm.sv"
`include "../env/svbt_data_in_generator.sv"
`include "../env/svbt_data_in_bfm.sv"
`include "../env/svbt_channel_out_generator.sv"
`include "../env/svbt_channel_out_bfm.sv"
`include "../env/svbt_environment.sv"

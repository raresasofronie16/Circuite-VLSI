
`include "svbt_interface.sv"
`include "svbt_base_unit.sv"
`include "svbt_packet.sv"
`include "svbt_reset_bfm.sv"
`include "svbt_data_in_generator.sv"
`include "svbt_data_in_bfm.sv"
`include "svbt_channel_out_generator.sv"
`include "svbt_channel_out_bfm.sv"
`include "svbt_environment.sv"

`include "router.v"

module top_inst(clock, reset, packet_valid, data, channel0, channel1, channel2, vld_chan_0, vld_chan_1, vld_chan_2, read_enb_0, read_enb_1, read_enb_2, suspend_data_in, err);
   input          clock;
   input          reset;
   input          packet_valid;
   input    [7:0] data;
   output   [7:0] channel0;
   output   [7:0] channel1;
   output   [7:0] channel2;
   output         vld_chan_0;
   output         vld_chan_1;
   output         vld_chan_2;
   input          read_enb_0;
   input          read_enb_1;
   input          read_enb_2;
   output         suspend_data_in;
   output         err;

   router router1 (.clk             (clock), // input
                   .reset_b         (reset), // input
                   .packet_valid    (packet_valid), // input
                   .data            (data), // input
                   .channel0        (channel0), // output
                   .vld_chan_0      (vld_chan_0), // output
                   .read_enb_0      (read_enb_0), // input
                   
                   //LAB: Tie together the signals for output interfaces 1 and 2
                   //(hint: look in hdl/router.v to see the signals declared in the top design file)
                   .channel1(channel1),
                   .vld_chan_1(vld_chan_1),
                   .read_enb_1(read_enb_1),
                   
                   .channel2(channel2),
                   .vld_chan_2(vld_chan_2),
                   .read_enb_2(read_enb_2),
                   
                   .suspend_data_in (suspend_data_in), // output
                   .err             (err)); // output

   reset_intf reset_intf(
      .clock(clock),
      .reset(reset)
   );
   
   input_intf input_intf(
      .clock(clock),
      .packet_valid(packet_valid),
      //LAB: Add the rest of the signals for this interface
     .data(data),
     .err(err),
     .suspend_data_in(suspend_data_in)
   );
   
   output_intf output_intf0(
      .clock(clock),
      .channel(channel0),
      .vld_chan(vld_chan_0),
      .read_enb(read_enb_0)
   );

  //LAB: Instantiate the rest of the output interfaces
     output_intf output_intf1(
      .clock(clock),
       .channel(channel1),
       .vld_chan(vld_chan_1),
       .read_enb(read_enb_1)
   );
     output_intf output_intf2(
      .clock(clock),
       .channel(channel2),
       .vld_chan(vld_chan_2),
       .read_enb(read_enb_2)
   );


endmodule

`include "../env/svbt_interface.sv"
`include "../env/svbt_base_unit.sv"
`include "../env/svbt_packet.sv"
`include "../env/svbt_environment.sv"

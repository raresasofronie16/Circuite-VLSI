// // Code your design here
// `include "svbt_interface.sv"
// `include "svbt_packet.sv"